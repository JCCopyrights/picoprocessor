-----------------------------------------------------------------------------
-- @(#) File: pico_types.vhd                                               --
-----------------------------------------------------------------------------
-- Authors: Yago Torroja                                yago@etsii.upm.es  --
-----------------------------------------------------------------------------
-- Copyright Universidad Politecnica de Madrid                             --
-----------------------------------------------------------------------------
-- E.T.S. de Ingenieros Industriales                                       --
-- Division de Ingenieria Electronica (UPM-DIE)                            --
-- E.T.S.I Industriales                                                    --
-- Jose Gutierrez Abascal, 2                                               --
-- MADRID 28006                                                            --
-- Tel : +34-1-3363191/92/93/94   Fax : +34-1-5645966                      --
-----------------------------------------------------------------------------
-- PROJECT: picoProcessor                                                  --
--                                                                         --
-----------------------------------------------------------------------------
-- Block      |                                                            --
--            |                                                            --
-- Description| BASIC TYPES                                                --
--            |                                                            --
-- Parameters |                                                            --
--            |                                                            --
-----------------------------------------------------------------------------
-- Dependencies:                                                           --
--               std_logic_1164                                            --
--                                                                         --
-----------------------------------------------------------------------------
-- Comments:                                                               --
--                                                                         --
-----------------------------------------------------------------------------
-- Version: 1.0                                        Fecha:              --
-----------------------------------------------------------------------------
-- Ver  |  Date    | Auth  | Version description                           --
--------|----------|-------|-------------------------------------------------
--      | 28/02/05 |  YT   | FIRST VERSION                                 --
--      |          |       |                                               --
-----------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

package pico_types is

----------------------------------------------------------------------------
-- General definitions, constants and types
----------------------------------------------------------------------------
  constant  AddrWidth   : natural := 12;
  constant  DataWidth   : natural := 8;

end pico_types;










